module PATTERN_Decoder3x8 (
    input [2:0] address,
    output [7:0] pattern
);
    
endmodule