`include "PATTERN_Decoder3x8.v"
`include "Decoder3x8.v"
module TESTBED ();
    
endmodule