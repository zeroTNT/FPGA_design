// File: PATTERN_Decoder3x8.v
// Generated with: v1.0.0
// Last update: 2025-02-20 21:09
//###########################################################################
// Design unit: PATTERN_Decoder3x8
//###########################################################################
// Purpose: This module is a 3x8 decoder that generates a pattern based on the input address.
//###########################################################################

module PATTERN_Decoder3x8 (
    input [2:0] address,
    output [7:0] pattern
);
    
endmodule