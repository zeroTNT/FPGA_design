// File: TESTBED.v
// Generated with: v1.0.0
// Last update: 2025-02-20 21:09
//###########################################################################
// Design unit: TESTBED
//###########################################################################
// Purpose: This module is a test bench for the PATTERN_Decoder3x8 module.
//###########################################################################
`include "PATTERN_Decoder3x8.v"
`include "Decoder3x8.v"
module TESTBED ();
    
endmodule